`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   11:08:43 03/11/2018
// Design Name:   f_alu
// Module Name:   /home/ise/Desktop/kek/fp_alu/falu_tb.v
// Project Name:  fp_alu
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: f_alu
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module falu_tb;

	// Inputs
	reg [31:0] a,b,a1,b1;
	reg clk,f;
	reg [2:0] op,op1;
	// Outputs
	wire [31:0] out;

	// Instantiate the Unit Under Test (UUT)
	float_alu uut (
		.a(a),.b(b),.clk(clk),.op(op), 
		.out(out)
	);
	always #5 clk=~clk;
	
	always@(posedge clk) begin
		a1<=repeat(2) @(posedge clk) a;
		b1<=repeat(2) @(posedge clk)b;
		op1<=repeat(2) @(posedge clk)op;
	end
	
	always@(posedge clk)
		$display("op=%b,a=%b %b %b,b=%b %b %b,c=%b %b %b",op1,a1[31],a1[30:23],a1[22:0],b1[31],b1[30:23],b1[22:0],out[31],out[30:23],out[22:0]);
	
	initial begin
		// Initialize Inputs
		clk=0;f=0;
		
		b=32'b0_10000000_00000000000000000000000;
		
		op=0;
		a=32'b0_10000001_11010000000000000000000;
		#10;
		a=32'b0_01111011_11010000000000000000000;
		#10;
		a=32'b0_01111111_11010000000000000000000;
		#50;	
		
		op=1;
		a=32'b0_10000001_11010000000000000000000;
		#10;
		a=32'b0_01111011_11010000000000000000000;
		#10;
		a=32'b0_01111111_11010000000000000000000;
		#50;
		
		op=2;
		a=32'b0_10000001_11010000000000000000000;
		#10;
		a=32'b0_01111011_11010000000000000000000;
		#10;
		a=32'b0_01111111_11010000000000000000000;
		#50;
		
		op=3;
		a=32'b0_10000001_11010000000000000000000;
		#10;
		a=32'b0_01111011_11010000000000000000000;
		#10;
		a=32'b0_01111111_11010000000000000000000;
		#50;
		
		op=4;
		a=32'b0_10000001_11010000000000000000000;
		#10;
		a=32'b0_01111011_11010000000000000000000;
		#10;
		a=32'b0_01111111_11010000000000000000000;
		#50;
		
		op=5;
		a=32'b0_10000001_11010000000000000000000;
		#10;
		a=32'b0_01111011_11010000000000000000000;
		#10;
		a=32'b0_01111111_11010000000000000000000;
		#50;
		
		op=6;
		a=32'b0_10000001_11010000000000000000000;
		#10;
		a=32'b0_01111011_11010000000000000000000;
		#10;
		a=32'b0_01111111_11010000000000000000000;
		#50;
		
		op=7;
		a=32'b0_10000001_11010000000000000000000;
		#10;
		a=32'b0_01111011_11010000000000000000000;
		#10;
		a=32'b0_01111111_11010000000000000000000;
		#50;
		
		$finish;
	end
      
endmodule

